`include "network_parms.h"
module mult_adder(
      input     clock, 
		  input     reset, 
		  input [`MULT_ADDER_IN_BITWIDTH:0]  in,
		  input [`MULT_ADDER_IN_BITWIDTH:0]  kernal,
		  output [`CONV_PRODUCT_WIDTH:0] out	
		  );

// wire declarations
wire [`CONV_PRODUCT_WIDTH:0] in_add_vector_wire [`KERNEL_SIZE_SQ];
wire [`CONV_PRODUCT_WIDTH:0] adder_tree_wire [(`KERNEL_SIZE_SQ*2)-1];
wire carry_wire [(`KERNEL_SIZE_SQ*2)-1];  

// assign statments
assign out = adder_tree_wire[0];
assign carry_wire [(`KERNEL_SIZE_SQ*2)-1-1:`KERNEL_SIZE_SQ-1] = `KERNEL_SIZE_SQ'd0;

// connect input vector to multipliers
genvar i;
generate
for(i = 0; i < `KERNEL_SIZE_SQ; i=i+1) begin : connect_mul
   mult_adder_mult ma_mult_inst(
    .clock(clock),
    .reset(reset),
    .operand_a([`CONV_MULT_WIDTH*(i+1)-1:i*`CONV_MULT_WIDTH]in),
    .operand_b([`CONV_MULT_WIDTH*(i+1)-1:i*`CONV_MULT_WIDTH]kernal),
    .out(in_add_vector_wire[i])
			     ); 
  end
endgenerate

// map products to adder tree wire
genvar i;
generate
for(i = 0; i < `KERNEL_SIZE_SQ; i=i+1) begin : connect_in_vector
    assign adder_tree_wire[i+`KERNEL_SIZE_SQ-1] = { `MA_ADDER_TREE_PAD'd0,
      in[(`CONV_PRODUCT_WIDTH*i)+`CONV_PRODUCT_BITWIDTH:`CONV_PRODUCT_WIDTH*i] };
  end
endgenerate

// connect adder tree
genvar j;
generate
for(j= (`KERNIL_SIZE_SQ*2)-2 ; j >=1 ; j=j-2) begin : sum_products
  mult_adder_add ma_add_inst(
    .clock(clock),
    .reset(reset),
    .operand_a(adder_tree_wire[j-1]),
    .operand_b(adder_tree_wire[j]),
    .c_a(carry_wire[j-1]),
    .c_b(carry_wire[j]),
    .out(adder_tree_wire[(j/2)-1]),
    .carry(carry_wire[(j/2)-1])
  );  

end // for
endgenerate
   
endmodule // mult_adder

module mult_adder_mult(
  input clock,
  input reset,
  input [`CONV_MULT_WIDTH:0] operand_a,
  input [`CONV_MULT_WIDTH:0] operand_b,
  output [`CONV_PRODUCT_WIDTH:0] out 
);
   reg [`CONV_PRODUCT_WIDTH:0]    product;
   
   assign out = product[`CONV_PRODUCT_WIDTH:0];

   always@(posedge clock or negedge reset) begin
      if(reset == 1'b0) 
	      product <= `CONV_PRODUCT_WIDTH'd0;
      else  
	      product <= operand_a * operand_b;
   end // always
endmodule

module mult_adder_add(
  input clock,
  input reset,
  input [`CONV_PRODUCT_WIDTH:0] operand_a,
  input [`CONV_PRODUCT_WIDTH:0] operand_b,
  input c_a, // overflow or carry indicators
  input c_b,
  output [`CONV_PRODUCT_WIDTH:0] out,
  output carry
);
   reg [`CONV_PRODUCT_WIDTH+1:0]    sum;

   assign out = sum[`CONV_PRODUCT_WIDTH:0];
   assign carry = sum[`CONV_PRODUCT_WIDTH+1] | c_a | c_b;
   
   always@(posedge clock or negedge reset) begin
      if(reset == 1'b0) 
	      sum <= `CONV_MULT_WIDTH'd0;
      else  
	      sum <= operand_a + operand_b;
   end // always
   endmodule
