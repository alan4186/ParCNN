module bus
(
  clk,
  rst,
  en, // an enable signal to start feeding data to FFT
  rom_data,
  rom_addr,
  pOut,
  nextSampleBtn,
  full_row
);
parameter bitWidth = 16,
          bw = bitWidth - 1,
          im_size = 28,
          im_s = im_size -1,
          rom_addr_size = 32; // needs to be changed!!!!!!!!!!

integer i,j,k;

input clk, rst, en, nextSampleBtn;
input [bw:0] rom_data;
input [1 + 9:0] rom_addr;

output full_row;
output [bw:0] pOut [0:im_s];

reg [4:0] row_count;
reg [bw:0] pOut [0:im_s];
reg [bw:0] test_reg [0:im_s];

always@(posedge clk or negedge rst) begin
  if(rst == 1'b0) begin
    for(i=0;i<im_size;i=i+1) begin
      pOut <= bw'd0;
    end
    rom_addr <= rom_addr_size'd0;
    ss <= 4'd0;
    full_row <= 1'b0;
  ////////////////////////////////////////
  //        next sample button
  ////////////////////////////////////////
  end else if (nextSampleBtn == 1'b1) begin
    rom_addr <= rom_addr_size'd0; 
    ss <= ss + 4'd1;
  ////////////////////////////////////////
  //      shift in data
  ////////////////////////////////////////
  end else if(read_rom == 1'b1) begin
    if(row_count <= 5'd28) begin
      pOut[0] <= rom_data;
      for(j=1;j<im_size;j=j+1) begin
        pOut[j] <= pOut[j-1]; // shift
      end
      rom_addr <= rom_addr + rom_addr_size'd1;
      row_count <= row_count + 5'd1;
      full_row <= 1'b0;
    end else begin
      row_count <= 5'd0;
      full_row <= 1'b1;
      for(k=0;k<im_size;k=k+1) begin
        test_reg[k] <= pOut[k];
      end
    end
  end
    
end
endmodule
